module D_ff ( 
    input  wire clk, rst, D, 
    output reg  Q 
); 
    always @(posedge clk or posedge rst) begin 
        if (rst) 
            Q <= 1'b0;   // Reset 
        else 
            Q <= D;      // Capture D at clock edge 
    end 
endmodule